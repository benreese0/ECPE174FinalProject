/***************************************************************
 * Game Logic
 * 
 * This top level files brings all the pong files together and 
 * runs the actual game.
 * 
 * Project: ECPE 174: Advanced Digital Design Final Project
 * Author:Jennifer Valencia
 * Date: 2013-11-08
 ***************************************************************/