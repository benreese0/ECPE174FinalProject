/***************************************************************
 * Paddle
 * 
 * <DESCRIPTION OF FILE>
 * 
 * Project: ECPE 174: Advanced Digital Design Final Project
 * Author:<AUTHOR NAME>
 * Date: 2013-11-08
 ***************************************************************/