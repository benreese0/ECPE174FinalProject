/***************************************************************
 * Audio
 * 
 * Sends output to WM8731
 * 
 * Project: ECPE 174: Advanced Digital Design Final Project
 * Author:Ben Reese
 * Date: 2013-11-08
 ***************************************************************/
 
 module Audio(input logic wall_hit, paddle_hit, point, win ,
				input logic lvl_up, clk,
				output logic m_clock);
/*				
audioclockdiv m_clock_gen(.iclk(clk), .oclk(m_clcok));
AUD_ADCLRCK
AUD_ADCDAT
AUD_DACLRCK
AUD_DACDAT
AUD_XCK
AUD_BCLK
I2C_SCLK
I2C_SDAT*/
				
				
endmodule
