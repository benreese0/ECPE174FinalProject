/***************************************************************
 * Constants
 * 
 * Has project wide constants defined
 * 
 * Project: ECPE 174: Advanced Digital Design Final Project
 * Author:Ben Reese
 * Date: 2013-11-08
 ***************************************************************/
 
 //Using sxample SVGA resolution
 const int X_RESOLUTION = 800;
 const int Y_RESOLUTION = 600;
 
 //Don't want the paddle to go cray-cray
 //~1/4 second to go from bottom to top of screen
 const int PADDLE_TICKS_PER_PIXEL = 20000;
 