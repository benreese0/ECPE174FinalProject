/***************************************************************
 * Ball
 * 
 * The following file tracks the ball position, the integer output
 * is the center pixel of the ball.
 * 
 * Project: ECPE 174: Advanced Digital Design Final Project
 * Author:Jennifer Valencia 
 * Date: 2013-11-08
 ***************************************************************/
 module Ball(input logic clk, rst);
 
 always_ff @ (posedge clk or negedge rst) begin
 
 
 endmodule
 